module inverse_table
#(parameter DIVISOR_WIDTH=7,WIDTH_INVERSE=8,WIDTH_SHIFT=4)
(
input [ DIVISOR_WIDTH-1:0] divisor,

output reg [WIDTH_INVERSE-1:0] div_inverse,
output reg [  WIDTH_SHIFT-1:0] div_shift
);

//inverses here all have 8 effective bits (the leftmost bit is 1)
always@* begin
	case(divisor)
	  7'd1   : div_inverse = 8'd128;
	  7'd2   : div_inverse = 8'd128;
	  7'd3   : div_inverse = 8'd171;
	  7'd4   : div_inverse = 8'd128;
	  7'd5   : div_inverse = 8'd205;
	  7'd6   : div_inverse = 8'd171;
	  7'd7   : div_inverse = 8'd147;
	  7'd8   : div_inverse = 8'd128;
	  7'd9   : div_inverse = 8'd228;
	  7'd10  : div_inverse = 8'd205;
	  7'd11  : div_inverse = 8'd187;
	  7'd12  : div_inverse = 8'd171;
	  7'd13  : div_inverse = 8'd158;
	  7'd14  : div_inverse = 8'd147;
	  7'd15  : div_inverse = 8'd137;
	  7'd16  : div_inverse = 8'd128;
	  7'd17  : div_inverse = 8'd241;
	  7'd18  : div_inverse = 8'd228;
	  7'd19  : div_inverse = 8'd216;
	  7'd20  : div_inverse = 8'd205;
	  7'd21  : div_inverse = 8'd196;
	  7'd22  : div_inverse = 8'd187;
	  7'd23  : div_inverse = 8'd179;
	  7'd24  : div_inverse = 8'd171;
	  7'd25  : div_inverse = 8'd164;
	  7'd26  : div_inverse = 8'd158;
	  7'd27  : div_inverse = 8'd152;
	  7'd28  : div_inverse = 8'd147;
	  7'd29  : div_inverse = 8'd142;
	  7'd30  : div_inverse = 8'd137;
	  7'd31  : div_inverse = 8'd133;
	  7'd32  : div_inverse = 8'd128;
	  7'd33  : div_inverse = 8'd249;
	  7'd34  : div_inverse = 8'd241;
	  7'd35  : div_inverse = 8'd235;
	  7'd36  : div_inverse = 8'd228;
	  7'd37  : div_inverse = 8'd222;
	  7'd38  : div_inverse = 8'd216;
	  7'd39  : div_inverse = 8'd211;
	  7'd40  : div_inverse = 8'd205;
	  7'd41  : div_inverse = 8'd200;
	  7'd42  : div_inverse = 8'd196;
	  7'd43  : div_inverse = 8'd191;
	  7'd44  : div_inverse = 8'd187;
	  7'd45  : div_inverse = 8'd183;
	  7'd46  : div_inverse = 8'd179;
	  7'd47  : div_inverse = 8'd175;
	  7'd48  : div_inverse = 8'd171;
	  7'd49  : div_inverse = 8'd168;
	  7'd50  : div_inverse = 8'd164;
	  7'd51  : div_inverse = 8'd161;
	  7'd52  : div_inverse = 8'd158;
	  7'd53  : div_inverse = 8'd155;
	  7'd54  : div_inverse = 8'd152;
	  7'd55  : div_inverse = 8'd149;
	  7'd56  : div_inverse = 8'd147;
	  7'd57  : div_inverse = 8'd144;
	  7'd58  : div_inverse = 8'd142;
	  7'd59  : div_inverse = 8'd139;
	  7'd60  : div_inverse = 8'd137;
	  7'd61  : div_inverse = 8'd135;
	  7'd62  : div_inverse = 8'd133;
	  7'd63  : div_inverse = 8'd131;
	  7'd64  : div_inverse = 8'd128;
	  7'd65  : div_inverse = 8'd253;
	  7'd66  : div_inverse = 8'd249;
	  7'd67  : div_inverse = 8'd245;
	  7'd68  : div_inverse = 8'd241;
	  7'd69  : div_inverse = 8'd238;
	  7'd70  : div_inverse = 8'd235;
	  7'd71  : div_inverse = 8'd231;
	  7'd72  : div_inverse = 8'd228;
	  7'd73  : div_inverse = 8'd225;
	  7'd74  : div_inverse = 8'd222;
	  7'd75  : div_inverse = 8'd219;
	  7'd76  : div_inverse = 8'd216;
	  7'd77  : div_inverse = 8'd213;
	  7'd78  : div_inverse = 8'd211;
	  7'd79  : div_inverse = 8'd208;
	  7'd80  : div_inverse = 8'd205;
	  7'd81  : div_inverse = 8'd203;
	  7'd82  : div_inverse = 8'd200;
	  7'd83  : div_inverse = 8'd198;
	  7'd84  : div_inverse = 8'd196;
	  7'd85  : div_inverse = 8'd193;
	  7'd86  : div_inverse = 8'd191;
	  7'd87  : div_inverse = 8'd189;
	  7'd88  : div_inverse = 8'd187;
	  7'd89  : div_inverse = 8'd185;
	  7'd90  : div_inverse = 8'd183;
	  7'd91  : div_inverse = 8'd181;
	  7'd92  : div_inverse = 8'd179;
	  7'd93  : div_inverse = 8'd177;
	  7'd94  : div_inverse = 8'd175;
	  7'd95  : div_inverse = 8'd173;
	  7'd96  : div_inverse = 8'd171;
	  7'd97  : div_inverse = 8'd169;
	  7'd98  : div_inverse = 8'd168;
	  7'd99  : div_inverse = 8'd166;
	  7'd100 : div_inverse = 8'd164;
	  7'd101 : div_inverse = 8'd163;
	  7'd102 : div_inverse = 8'd161;
	  7'd103 : div_inverse = 8'd160;
	  7'd104 : div_inverse = 8'd158;
	  7'd105 : div_inverse = 8'd157;
	default : div_inverse = 8'd128 ;  
  endcase
end


always@* begin
	case(divisor)
	  7'd1   : div_shift = 4'd7 ;
	  7'd2   : div_shift = 4'd8 ;
	  7'd3   : div_shift = 4'd9 ;
	  7'd4   : div_shift = 4'd9 ;
	  7'd5   : div_shift = 4'd10;
	  7'd6   : div_shift = 4'd10;
	  7'd7   : div_shift = 4'd10;
	  7'd8   : div_shift = 4'd10;
	  7'd9   : div_shift = 4'd11;
	  7'd10  : div_shift = 4'd11;
	  7'd11  : div_shift = 4'd11;
	  7'd12  : div_shift = 4'd11;
	  7'd13  : div_shift = 4'd11;
	  7'd14  : div_shift = 4'd11;
	  7'd15  : div_shift = 4'd11;
	  7'd16  : div_shift = 4'd11;
	  7'd17  : div_shift = 4'd12;
	  7'd18  : div_shift = 4'd12;
	  7'd19  : div_shift = 4'd12;
	  7'd20  : div_shift = 4'd12;
	  7'd21  : div_shift = 4'd12;
	  7'd22  : div_shift = 4'd12;
	  7'd23  : div_shift = 4'd12;
	  7'd24  : div_shift = 4'd12;
	  7'd25  : div_shift = 4'd12;
	  7'd26  : div_shift = 4'd12;
	  7'd27  : div_shift = 4'd12;
	  7'd28  : div_shift = 4'd12;
	  7'd29  : div_shift = 4'd12;
	  7'd30  : div_shift = 4'd12;
	  7'd31  : div_shift = 4'd12;
	  7'd32  : div_shift = 4'd12;
	  7'd33  : div_shift = 4'd13;
	  7'd34  : div_shift = 4'd13;
	  7'd35  : div_shift = 4'd13;
	  7'd36  : div_shift = 4'd13;
	  7'd37  : div_shift = 4'd13;
	  7'd38  : div_shift = 4'd13;
	  7'd39  : div_shift = 4'd13;
	  7'd40  : div_shift = 4'd13;
	  7'd41  : div_shift = 4'd13;
	  7'd42  : div_shift = 4'd13;
	  7'd43  : div_shift = 4'd13;
	  7'd44  : div_shift = 4'd13;
	  7'd45  : div_shift = 4'd13;
	  7'd46  : div_shift = 4'd13;
	  7'd47  : div_shift = 4'd13;
	  7'd48  : div_shift = 4'd13;
	  7'd49  : div_shift = 4'd13;
	  7'd50  : div_shift = 4'd13;
	  7'd51  : div_shift = 4'd13;
	  7'd52  : div_shift = 4'd13;
	  7'd53  : div_shift = 4'd13;
	  7'd54  : div_shift = 4'd13;
	  7'd55  : div_shift = 4'd13;
	  7'd56  : div_shift = 4'd13;
	  7'd57  : div_shift = 4'd13;
	  7'd58  : div_shift = 4'd13;
	  7'd59  : div_shift = 4'd13;
	  7'd60  : div_shift = 4'd13;
	  7'd61  : div_shift = 4'd13;
	  7'd62  : div_shift = 4'd13;
	  7'd63  : div_shift = 4'd13;
	  7'd64  : div_shift = 4'd13;
	  7'd65  : div_shift = 4'd14;
	  7'd66  : div_shift = 4'd14;
	  7'd67  : div_shift = 4'd14;
	  7'd68  : div_shift = 4'd14;
	  7'd69  : div_shift = 4'd14;
	  7'd70  : div_shift = 4'd14;
	  7'd71  : div_shift = 4'd14;
	  7'd72  : div_shift = 4'd14;
	  7'd73  : div_shift = 4'd14;
	  7'd74  : div_shift = 4'd14;
	  7'd75  : div_shift = 4'd14;
	  7'd76  : div_shift = 4'd14;
	  7'd77  : div_shift = 4'd14;
	  7'd78  : div_shift = 4'd14;
	  7'd79  : div_shift = 4'd14;
	  7'd80  : div_shift = 4'd14;
	  7'd81  : div_shift = 4'd14;
	  7'd82  : div_shift = 4'd14;
	  7'd83  : div_shift = 4'd14;
	  7'd84  : div_shift = 4'd14;
	  7'd85  : div_shift = 4'd14;
	  7'd86  : div_shift = 4'd14;
	  7'd87  : div_shift = 4'd14;
	  7'd88  : div_shift = 4'd14;
	  7'd89  : div_shift = 4'd14;
	  7'd90  : div_shift = 4'd14;
	  7'd91  : div_shift = 4'd14;
	  7'd92  : div_shift = 4'd14;
	  7'd93  : div_shift = 4'd14;
	  7'd94  : div_shift = 4'd14;
	  7'd95  : div_shift = 4'd14;
	  7'd96  : div_shift = 4'd14;
	  7'd97  : div_shift = 4'd14;
	  7'd98  : div_shift = 4'd14;
	  7'd99  : div_shift = 4'd14;
	  7'd100 : div_shift = 4'd14;
	  7'd101 : div_shift = 4'd14;
	  7'd102 : div_shift = 4'd14;
	  7'd103 : div_shift = 4'd14;
	  7'd104 : div_shift = 4'd14;
	  7'd105 : div_shift = 4'd14;
	default : div_shift = 4'd7 ;  
  endcase
end

endmodule